// AES Module
// This module implements an AES encryption and decryption system.
// It includes key expansion, encryption, and decryption stages.

module AES (
    input wire clk,                  // Clock signal
    input wire reset,                // Active-high reset signal
    input wire enable,               // Enable signal for encryption
    input wire [127:0] key128,       // 128-bit AES encryption key
    input wire [127:0] data_in,      // 128-bit data input (plaintext)

    output wire [127:0] encrypted_out, // 128-bit encrypted data output (ciphertext)
    output wire [127:0] decrypted_out  // 128-bit decrypted data output (plaintext)
);

    // Internal signals

    // aesReset128: Internal reset signal derived from the reset input
    wire aesReset128;

    // tempEncryptedOutput128: Temporary output wire for encrypted data from the AES encryption module
    wire [127:0] tempEncryptedOutput128;

    // tempDecryptedOutput128: Temporary output wire for decrypted data from the AES decryption module
    wire [127:0] tempDecryptedOutput128;

    // allKeys128: Wire holding the expanded keys generated by the KeyExpansion module
    // Size is 1408 bits for storing all round keys required by AES (128-bit key version)
    wire [1407:0] allKeys128;

    // Generate internal reset signal
    // This ensures aesReset128 is active when reset is active
    assign aesReset128 = reset;

    // Key Expansion Module for 128-bit AES
    // Generates expanded keys for encryption and decryption using the provided 128-bit key
    // Parameters (4, 10) specify AES with 4 columns and 10 rounds for 128-bit key
    KeyExpansion #(4, 10) keysGetter128 (
        .keyIn(key128),        // Input: original 128-bit key
        .keysOut(allKeys128)  // Output: all expanded round keys (1408 bits)
    );

    // AES Encryption Module
    // Encrypts the input data using the expanded keys
    // Parameters (4, 10) indicate 128-bit AES with 4 columns and 10 rounds
    AESEncrypt #(4, 10) aese128 (
        .data(data_in),             // Input: plaintext data to encrypt
        .allKeys(allKeys128),     // Input: expanded keys for encryption
        .state(tempEncryptedOutput128), // Output: encrypted data (ciphertext)
        .clk(clk),                     // Clock signal
        .enable(enable),               // Enable signal for encryption
        .reset(aesReset128)            // Reset signal
    );

    // AES Decryption Module
    // Decrypts the encrypted data to obtain the original plaintext
    // Parameters (4, 10) specify 128-bit AES with 4 columns and 10 rounds
    AESDecrypt #(4, 10) aesd128 (
        .data(tempEncryptedOutput128), // Input: encrypted data to decrypt (ciphertext)
        .allKeys(allKeys128),        // Input: expanded keys for decryption
        .state(tempDecryptedOutput128), // Output: decrypted data (plaintext)
        .clk(clk),                        // Clock signal
        .enable(enable),                  // Enable signal for decryption
        .reset(aesReset128)               // Reset signal
    );

    // Output assignments
    // Assigns the encrypted and decrypted data to the module outputs
    assign encrypted_out = tempEncryptedOutput128; // Encrypted data output
    assign decrypted_out = tempDecryptedOutput128; // Decrypted data output

endmodule
